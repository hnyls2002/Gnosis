module reorder_buffer(
    // cpu
    input wire  clk,
    input wire  rst,
    input wire  rdy

    // inst info
);
endmodule