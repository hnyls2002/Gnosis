module dispatcher(
);

endmodule