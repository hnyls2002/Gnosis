module decoder (
);
    
endmodule